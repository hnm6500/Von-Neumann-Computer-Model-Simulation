`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: 
// Engineer: 
// 
// Create Date:    16:43:14 02/20/2017 
// Design Name: 
// Module Name:    Registe_File 
// Project Name: 
// Target Devices: 
// Tool versions: 
// Description: 
//
// Dependencies: 
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Registe_File(
    input rd1,
    input rd2,
    input rst,
    input clk,
    input wr,
    input in,
    input we,
    output out1,
    output out2
    );


endmodule
